
module hx8352_controller_fsm(
	input clk,
	input rst,
	output init_done,
	output reg [15:0]data_to_write,
	output command_or_data,
	output bus_step,
	output wire [15:0]delay_value,
	output wire delay_step,
	output reg lcd_cs
);
localparam 
HIGH    = 1'b1,
LOW     = 1'b0,
LCD_CMD    = 1'b0,
LCD_DATA   = 1'b1,
CMD_Product_ID								=	8'h00,
CMD_Data_read_write						=	8'h22,
STATE_INITIALIZE							= 4'd1,
STATE_IDLE									= 4'd2,
STATE_TRANSFER_CMD 						= 4'd3,
STATE_TRANSFER_PIXEL						= 4'd4,
STATE_TRANSFER_PIXEL_LOAD_CMD 		= 4'd5,
STATE_TRANSFER_PIXEL_LOAD_CMD_END	= 4'd6,
STATE_TRANSFER_PIXEL_LOAD_DATA		= 4'd7,
STATE_TRANSFER_PIXEL_LOAD_DATA_END	= 4'd8

;


reg  lcd_init_step;
wire lcd_init_working;
wire lcd_bus_step;
wire lcd_command_or_data;
wire [15:0]lcd_data_to_write;
hx8352_lcd_init 
	init_ut0( 
	.clk(clk),
	.rst(rst),
	.step(lcd_init_step),
	.delay_step(delay_step),
	.delay_value(delay_value),
	.data_to_write(lcd_data_to_write),
	.command_or_data(lcd_command_or_data),
	.working(lcd_init_working),
	.done(init_done),
	.bus_step(lcd_bus_step)
	);
	
reg  [3:0]  fsm_state;
reg bus_step_reg;
reg command_or_data_reg;
always @(posedge clk or posedge rst) begin
  if (rst) begin
		fsm_state <= STATE_INITIALIZE;
		lcd_init_step <= LOW;
		data_to_write <= 16'h0000;
		bus_step_reg <= LOW;
		command_or_data_reg <= LCD_CMD;
		lcd_cs <= HIGH;
  end else begin 	
		lcd_init_step <= LOW;
		case (fsm_state)
			STATE_IDLE: begin
				//if(step_sync) begin
					//if(write_cmd_reg)
						//fsm_state <= STATE_TRANSFER_CMD;
					//else

				lcd_cs <= HIGH;
				fsm_state <= STATE_TRANSFER_PIXEL;
				//end
			end
			//STATE_TRANSFER_CMD: begin
			//	bus_step <= HIGH;
			//	case (pc)
			//		8'h00:  
			//		8'h01:  {pc,command_or_data, data_to_write}     <= {pc+1,LCD_CMD,  {8'h00, cmd_in_reg}}; 
			//		8'h02:  {pc,command_or_data, data_to_write}     <= {pc+1,LCD_DATA, data_in_reg}; 
			//		8'h03:  begin //! NOP
			//				command_or_data <= LCD_CMD;
			//				data_to_write <= {8'h00, CMD_Product_ID};
			//				fsm_state <= STATE_IDLE;						
			//				end
			//		default: fsm_state <= STATE_IDLE; 
			//	endcase
			//end			
			STATE_TRANSFER_PIXEL: begin
				bus_step_reg <= LOW;
				fsm_state <= STATE_IDLE; 
			end
			STATE_TRANSFER_PIXEL_LOAD_CMD : begin
				command_or_data_reg <= LCD_CMD;
				data_to_write   <= {8'h00, CMD_Data_read_write};
				bus_step_reg <= HIGH;
				fsm_state <= STATE_TRANSFER_PIXEL_LOAD_CMD_END; 
			end 
			STATE_TRANSFER_PIXEL_LOAD_CMD_END : begin
				bus_step_reg <= LOW;
				fsm_state <= STATE_TRANSFER_PIXEL_LOAD_DATA; 
			end
			STATE_TRANSFER_PIXEL_LOAD_DATA: begin 
				command_or_data_reg <= LCD_DATA;
				data_to_write <= {16'hAABB};
				bus_step_reg <= HIGH;
				fsm_state <= STATE_TRANSFER_PIXEL_LOAD_DATA_END; 
			end
			STATE_TRANSFER_PIXEL_LOAD_DATA_END : begin
				command_or_data_reg <= LCD_CMD;
				data_to_write <= {8'h00, CMD_Product_ID};
				bus_step_reg <= LOW;
				fsm_state <= STATE_IDLE; 
			end
			STATE_INITIALIZE: begin
				lcd_cs <= LOW;
				if(init_done)
					fsm_state <= STATE_IDLE;
				else if(!lcd_init_working) begin
					lcd_init_step <= 1'b1;
				end
				if(lcd_bus_step) begin
					data_to_write <= lcd_data_to_write;
					command_or_data_reg <= lcd_command_or_data;
				end
			end
		default: fsm_state <= STATE_INITIALIZE;
		endcase
	end
end
 
assign bus_step = lcd_bus_step | bus_step_reg;
assign command_or_data = command_or_data_reg;
endmodule 


module hx8352_lcd_init( 
	input  clk,
	input  rst,
	input  step,
	output reg delay_step,
	output reg [15:0]delay_value,
	output reg command_or_data,
	output reg [15:0]data_to_write,
	output working,
	output done,
	output bus_step
	);
localparam 
HIGH    = 1'b1,
LOW     = 1'b0,
LCD_CMD    = 1'b0,
LCD_DATA   = 1'b1,
/* 6.1 Command set = Taken from datasheet */
CMD_Product_ID								=	8'h00,
CMD_Display_mode							=	8'h01,
CMD_Column_Address_Start_1				=	8'h02,
CMD_Column_Address_Start_2				=	8'h03,
CMD_Column_Address_End_1				=	8'h04,
CMD_Column_Address_End_2				=	8'h05,
CMD_Row_Address_Start_1					=	8'h06,
CMD_Row_Address_Start_2					=	8'h07,
CMD_Row_Address_End_1					=	8'h08,
CMD_Row_Address_End_2					=	8'h09,
CMD_Partial_Area_Start_Row_1			=	8'h0a,
CMD_Partial_Area_Start_Row_2			=	8'h0b,
CMD_Partial_Area_End_Row_1				=	8'h0c,
CMD_Partial_Area_End_Row_2				=	8'h0d,
CMD_Vertical_Scroll_Top_Fixed_Area_1=	8'h0e,
CMD_Vertical_Scroll_Top_Fixed_Area_2=	8'h0f,
CMD_Vertical_Scroll_Height_Area_1	=	8'h10,
CMD_Vertical_Scroll_Height_Area_2	=	8'h11,
CMD_Vertical_Scroll_Button_Fixed_1	=	8'h12,
CMD_Vertical_Scroll_Button_Fixed_2	=	8'h13,
CMD_Vertical_Scroll_Start_Address_1	=	8'h14,
CMD_Vertical_Scroll_Start_Address_2	=	8'h15,
CMD_Memory_Access_Control				=	8'h16,
CMD_OSC_Control_1							=	8'h17,
CMD_OSC_Control_2							=	8'h18,
CMD_Power_Control_1						=	8'h19,
CMD_Power_Control_2						=	8'h1a,
CMD_Power_Control_3						=	8'h1b,
CMD_Power_Control_4						=	8'h1c,
CMD_Power_Control_5						=	8'h1d,
CMD_Power_Control_6						=	8'h1e,
CMD_VCOM_Control							=	8'h1f,
CMD_Data_read_write						=	8'h22,
CMD_Display_Control_1					=	8'h23,
CMD_Display_Control_2					=	8'h24,
CMD_Display_Control_3					=	8'h25,
CMD_Display_Control_4					=	8'h26,
CMD_Display_Control_5					=	8'h27,
CMD_Display_Control_6					=	8'h28,
CMD_Display_Control_7					=	8'h29,
CMD_Display_Control_8					=	8'h2a,
CMD_Cycle_Control_1						=	8'h2b,
CMD_Cycle_Control_2						=	8'h2c,
CMD_Cycle_Control_3						=	8'h2d,
CMD_Cycle_Control_4						=	8'h2e,
CMD_Cycle_Control_5						=	8'h2f,
CMD_Cycle_Control_6						=	8'h30,
CMD_Cycle_Control_7						=	8'h31,
CMD_Cycle_Control_8						=	8'h32,
CMD_Cycle_Control_10						=	8'h34,
CMD_Cycle_Control_11						=	8'h35,
CMD_Cycle_Control_12						=	8'h36,
CMD_Cycle_Control_13						=	8'h37,
CMD_Cycle_Control_14						=	8'h38,
CMD_Cycle_Control_15						=	8'h39,
CMD_Interface_Control_1					=	8'h3a,
CMD_Source_Control_1						=	8'h3c,
CMD_Source_Control_2						=	8'h3d,
CMD_Gamma_Control_1						=	8'h3e,
CMD_Gamma_Control_2						=	8'h3f,
CMD_Gamma_Control_3						=	8'h40,
CMD_Gamma_Control_4						=	8'h41,
CMD_Gamma_Control_5						=	8'h42,
CMD_Gamma_Control_6						=	8'h43,
CMD_Gamma_Control_7						=	8'h44,
CMD_Gamma_Control_8						=	8'h45,
CMD_Gamma_Control_9						=	8'h46,
CMD_Gamma_Control_10						=	8'h47,
CMD_Gamma_Control_11						=	8'h48,
CMD_Gamma_Control_12						=	8'h49,
CMD_PANEL_Control							=	8'h55,
CMD_OTP_1									=	8'h56,
CMD_OTP_2									=	8'h57,
CMD_OTP_3									=	8'h58,
CMD_OTP_4									=	8'h59,
CMD_IP_Control								=	8'h5a,
CMD_DGC_LUT_WRITE							=	8'h5c,
CMD_DATA_Control							=	8'h5d,
CMD_Test_Mode								=	8'h83,
CMD_VDDD_control							=	8'h85,
CMD_Powr_driving_Control				=	8'h8A,
CMD_VGS_RES_control_1					=	8'h8B,
CMD_VGS_RES_control_2					=	8'h8C,
CMD_PWM_Control_0							=	8'h91,
CMD_PWM_Control_1							=	8'h95,
CMD_PWM_Control_2							=	8'h96,
CMD_PWM_Control_3							=	8'h97,
CMD_CABC_Period_Control_1				=	8'h6B,
CMD_CABC_Period_Control_2				=	8'h6C,
CMD_CABC_Gain1								=	8'h6F,
CMD_CABC_Gain2								=	8'h70,
CMD_CABC_Gain3								=	8'h71,
CMD_CABC_Gain4								=	8'h72,
CMD_CABC_Gain5								=	8'h73,
CMD_CABC_Gain6								=	8'h74,
CMD_CABC_Gain7								=	8'h75,
CMD_CABC_Gain8								=	8'h76,
CMD_CABC_Gain9								=	8'h77,
PC_INDEX_DELAY_1							=	8'h4d,
PC_INDEX_DELAY_2							=	8'h5f,
PC_INDEX_DELAY_3							=	8'h69,
PC_INDEX_DELAY_4							=	8'h6f,
PC_INDEX_DELAY_5							=	8'h75,
PC_INDEX_DELAY_6							=	8'h8b,
PC_INDEX_DONE								=  8'hbd;

reg  [7:0] pc;
wire [7:0] pc_next;
reg enable;

always @(posedge clk or posedge rst) begin
	if (rst) begin
		enable <= 0;
	end
	else begin
		enable <= enable;
		if(step) 
			enable <= 1'b1;
		if(done) 
			enable <= 1'b0;
	end
end
wire enabled_clk;
assign enabled_clk = clk & enable; 
always @(posedge enabled_clk or posedge rst) begin
	if (rst) begin
		pc <= 0;
	end
	else begin
		pc <= pc_next;
	end
end

assign pc_next = (step) ? 1'b0 : pc + 1'b1;

always @(pc)
case (pc)
	8'h01:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Test_Mode}};
	8'h03:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h02}};//TESTM=1 
	8'h05:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_VDDD_control}};
	8'h07:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h03}};//VDC_SEL=011
	8'h09:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_VGS_RES_control_1}};
	8'h0b:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h01}};
	8'h0d:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_VGS_RES_control_2}};
	8'h0f:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h93}};//STBA[7]=1,STBA[5:4]=01,STBA[1:0]=11
	8'h11:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_PWM_Control_0}};
	8'h13:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h01}};//DCDC_SYNC=1
	8'h15:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Test_Mode}};
	8'h17:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h00}}; //TESTM=0

	8'h19:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Gamma_Control_1}};//Gamma Setting
	8'h1b:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'hB0}};
	8'h1d:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Gamma_Control_2}};
	8'h1f:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h03}};
	8'h21:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Gamma_Control_3}};
	8'h23:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h10}};
	8'h25:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Gamma_Control_5}};
	8'h27:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h13}};
	8'h29:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Gamma_Control_6}};
	8'h2b:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h46}};
	8'h2d:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Gamma_Control_7}};
	8'h2f:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h23}};
	8'h31:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Gamma_Control_8}};
	8'h33:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h76}};
	8'h35:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Gamma_Control_9}};
	8'h37:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h00}};
	8'h39:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Gamma_Control_10}};
	8'h3b:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h5E}};
	8'h3d:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Gamma_Control_11}};
	8'h3f:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h4F}};
	8'h41:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Gamma_Control_12}};
	8'h43:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h40}};

	8'h45:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00,CMD_OSC_Control_1}};//**********Power On sequence************
	8'h47:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h91}};
	8'h49:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Cycle_Control_1}};
	8'h4b:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'hF9}};
	PC_INDEX_DELAY_1:  
			  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'hF9}};//10ms delay
	8'h4f:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Power_Control_3}};
	8'h51:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h14}};
	8'h53:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Power_Control_2}};
	8'h55:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h11}};
	8'h57:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Power_Control_4}};
	8'h59:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h06}}; // 0d
	8'h5b:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_VCOM_Control}};
	8'h5d:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h42}};
	PC_INDEX_DELAY_2:  
			  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h42}};//20ms delay
	8'h61:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Power_Control_1}};
	8'h63:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h0A}};
	8'h65:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Power_Control_1}};
	8'h67:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h1A}};
	PC_INDEX_DELAY_3:  
			  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h1A}};//60ms delay
	8'h6a:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Power_Control_1}};
	8'h6c:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h12}};
	PC_INDEX_DELAY_4:  
	        {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h12}};//40ms delay
	8'h71:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Power_Control_6}};
	PC_INDEX_DELAY_5:  
			  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h27}};
	8'h75:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h27}};//60ms delay

	8'h77:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Display_Control_2}};//**********DISPLAY ON SETTING***********
	8'h79:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h60}};					
	8'h7b:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Source_Control_2}};
	8'h7d:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h40}};					
	8'h7f:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Cycle_Control_10}};
	8'h81:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h38}};					
	8'h83:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Cycle_Control_11}};
	8'h85:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h38}};					
	8'h87:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Display_Control_2}};
	8'h89:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h38}};
	PC_INDEX_DELAY_6:
			  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h38}};//40ms delay
	8'h8c:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Display_Control_2}};
	8'h8f:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h3C}};					
	8'h91:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Memory_Access_Control}};
	8'h93:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h1C}};					
	8'h95:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Display_mode}};
	8'h97:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h06}};					
	8'h99:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_PANEL_Control}};
	8'h9b:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h00}};					
	8'h9d:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Column_Address_Start_1}};
	8'h9f:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h00}};
	8'ha1:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Column_Address_Start_2}};
	8'ha3:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h00}};
	8'ha5:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Column_Address_End_1}};
	8'ha7:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h00}};
	8'ha9:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Column_Address_End_2}};
	8'hab:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'hEF}};					
	8'had:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Row_Address_Start_1}};
	8'haf:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h00}};
	8'hb1:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Row_Address_Start_2}};
	8'hb3:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h00}};
	8'hb5:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Row_Address_End_1}};
	8'hb7:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h01}};
	8'hb9:  {command_or_data, data_to_write}  = {LCD_CMD,  {8'h00, CMD_Row_Address_End_2}};
	8'hbb:  {command_or_data, data_to_write}  = {LCD_DATA, {8'h00, 8'h8F}};					
	8'hbd:  {command_or_data, data_to_write}  = {LCD_CMD, {8'h00, CMD_Product_ID}};  
	default: {command_or_data, data_to_write} = {LCD_CMD, 16'h0000}; 
endcase


always @(pc)
case (pc)
	PC_INDEX_DELAY_1: delay_value=15'd10_000;
	PC_INDEX_DELAY_2: delay_value=15'd20_000;
	PC_INDEX_DELAY_3: delay_value=15'd60_000;
	PC_INDEX_DELAY_4: delay_value=15'd40_000;
	PC_INDEX_DELAY_5: delay_value=15'd60_000;
	PC_INDEX_DELAY_6: delay_value=15'd40_000;
  default:delay_value=15'd0;
endcase
always @(pc)
case (pc)
	PC_INDEX_DELAY_1: delay_step=1'b1;
	PC_INDEX_DELAY_2: delay_step=1'b1;
	PC_INDEX_DELAY_3: delay_step=1'b1;
	PC_INDEX_DELAY_4: delay_step=1'b1;
	PC_INDEX_DELAY_5: delay_step=1'b1;
	PC_INDEX_DELAY_6: delay_step=1'b1;
  default:delay_step=1'b0;
endcase


assign done = pc == PC_INDEX_DONE;
assign working = enable;
assign bus_step = pc[0];

endmodule 